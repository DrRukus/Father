module main;
  initial
    begin
      $display("Goodbye, world!");
    end
endmodule
